----------------
--Problem 17.4--
----------------

